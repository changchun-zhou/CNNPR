module req2data_column_parallel #(
)
(
    input clk,
    input reset,
    input mode,
    input 
    output valid_index,
    )