library verilog;
use verilog.vl_types.all;
entity mem_controller_tb is
end mem_controller_tb;
